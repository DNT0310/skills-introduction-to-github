module helo;
endmodule
